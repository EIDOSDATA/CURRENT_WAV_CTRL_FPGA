`timescale 1ns/10ps


`define NOM_FREQ ("3.33")
	
/* Lattice XP2 internal Oscillator */	
/* NOM_FREQ: 2.08(default),2.15,2.22,2.29,2.38,2.46,2.56,2.66,2.77,2.89,
   3.02,3.17,3.33,3.50,3.69,3.91,4.16,4.29,4.43,4.59,4.75,4.93,5.12,5.32,5.54,
   5.78,6.05,6.33,6.65,7.00,7.39,7.82,8.31,8.58,8.87,9.17,9.50,9.85,10.23,10.64,
   11.08,11.57,12.09,12.67,13.30,14.00,14.78,15.65,16.63,17.73,19.00,20.46,
   22.17,24.18,26.60,29.56,33.25,38.00,44.33,53.20,66.50,88.67,133.00 MHz 
*/

module ci_stim_fpga_wrapper (	
	/**
	- FPGA related signals
	*/
	/* input ports */
	i_rst_n,
	//duty,
	
	/* output ports */		
	out_sw1_sig,
	out_sw2_sig,
	out_sw3_sig,
	out_sw4_sig,
	output_ctrl_sig	
) /* synthesis syn_force_pads=1 syn_noprune=1*/;
	/**
	- FPGA related signals
	*/
	/* input ports */
	input i_rst_n/* synthesis LOC="69" IO_TYPE="LVCMOS33" PULLMODE="UP" */;
	
	//input [7:0] duty/* synthesis LOC="25,24,21,20,19,18,17,16" IO_TYPE="LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33" PULLMODE="UP,UP,UP,UP,DOWN,DOWN,DOWN,DOWN" */; // 11110000
	//input [3:0] duty/* synthesis LOC="25,24,21,20" IO_TYPE="LVCMOS33,LVCMOS33,LVCMOS33,LVCMOS33" PULLMODE="DOWN,DOWN,UP,UP" */; // 0011
	
	/* output ports */	
	output out_sw1_sig/* synthesis LOC="64" IO_TYPE="LVCMOS33" PULLMODE="NONE" */; 
	output out_sw2_sig/* synthesis LOC="65" IO_TYPE="LVCMOS33" PULLMODE="NONE" */; 
	output out_sw3_sig/* synthesis LOC="66" IO_TYPE="LVCMOS33" PULLMODE="NONE" */;	
	output out_sw4_sig/* synthesis LOC="67" IO_TYPE="LVCMOS33" PULLMODE="NONE" */;
	output output_ctrl_sig/* synthesis LOC="68" IO_TYPE="LVCMOS33" PULLMODE="NONE" */;	
	
	reg out_sw1_sig;
	reg out_sw2_sig;
	reg out_sw3_sig;
	reg out_sw4_sig;
	reg output_ctrl_sig;
	/* internal wires and regs */
	/* IMPORTANT NOTES 
	  for specifying clock constraints, let SynplifyPro keep this wire name during synthesis by using this attribute
	*/
	wire w_clk 		/* synthesis syn_keep = 1 */;
	//wire w_div4_clk /* synthesis syn_keep = 1 */;
	//wire w_div64_clk 	/* synthesis syn_keep = 1 */;
	//wire w_div64x64_clk /* synthesis syn_keep = 1 */;
	//wire w_db_clk 	/* synthesis syn_keep = 1 */;
	//wire w_div64x4_clk /* synthesis syn_keep = 1 */;
	//wire w_slow_clk /* synthesis syn_keep = 1 */;
	
	/**
	- 1) Lattice IP instantiation
	    * Generates internal Clock and Reset
	*/
`ifdef SIMULATION
	/* Lattice GSR */
	//gsr GSR_INST (.gsr(i_rst_n));
		
	/* Lattice XP2 internal Oscillator */
	wire w_force_clk;

	assign w_clk = w_force_clk;
	//osch #(.NOM_FREQ(`NOM_FREQ))  internal_osc (.osc(w_clk));

`else
	/* Lattice GSR */
	/* GSR and PUR should make the instance name with pre-defined name which is "GSR_INST" and "PUR_INST" in each.
	   It is because their output is generated by Lattice tool and routed to all registers by the tool and so 
	   the tool should be able to find the instance automatically. This is the reason why instance name is fixed. */
	GSR GSR_INST (.GSR(i_rst_n));

//`define XO2

`ifdef XO2

	OSCH #(.NOM_FREQ(`NOM_FREQ))  internal_osc (.STDBY(1'b0), .OSC(w_clk), .SEDSTDBY());
`else

	/* Lattice XP2 internal Oscillator */	
	OSCE #(.NOM_FREQ(`NOM_FREQ))  internal_osc (.OSC(w_clk));
`endif
`endif
	
	reg [23:0] anode_duty = 3333; // 1ms
	reg [23:0] cathode_duty = 6999; // 3666 ~ 6999 >> 3333 >> 1ms
	reg [23:0] output_ctrl_duty = 6999; // +333
	reg [23:0] cnt_a;
	reg [23:0] cnt_c;
	reg [23:0] cnt_o;

    always @(posedge w_clk or negedge i_rst_n)
	begin
		if (~i_rst_n)begin
			cnt_a <= 0;
			cnt_c <= 0;
			cnt_o <= 0;
		end
		
		else if(cnt_a >= 3333333)begin //3333333 > 1sec
			cnt_a <= 0;
		end
		
		else if(cnt_c >= 3336999)begin //3336999 - 3666 = 3333333 >> 1sec
			cnt_c <= 3666; // anode after + 100us delay after
		end
		
		//else if(cnt_o >= 3336999)begin //3333333
			//cnt_o <= 3666;
		//end
		
		else begin
			cnt_a <= cnt_a + 1;
			cnt_c <= cnt_c + 1;
			cnt_o <= cnt_o + 1;
		end
	end
	
	// OUTPUT SW SIGNAL
	always @(posedge w_clk or negedge i_rst_n)
	begin
		if (~i_rst_n)begin
			out_sw1_sig <= 0;
			out_sw2_sig <= 0;
			out_sw3_sig <= 0;
			out_sw4_sig <= 0;			
		end
		
		else begin
			
			/* Anode SIGNAL */
			if(anode_duty >= cnt_a)begin
				out_sw1_sig <= 1;
				out_sw2_sig <= 1;				
			end
			else begin
				out_sw1_sig <= 0;
				out_sw2_sig <= 0;				
			end
			
			/* Cathode SIGNAL */
			if(cathode_duty >= cnt_c)begin
				out_sw3_sig <= 1;
				out_sw4_sig <= 1;				
			end
			else begin
				out_sw3_sig <= 0;
				out_sw4_sig <= 0;				
			end
			
			/* OUTPUT CTRL SIGNAL */
			if(3333 >= cnt_a || 6999 >= cnt_c)begin
				output_ctrl_sig <= 1;				
			end
			else begin
				output_ctrl_sig <= 0;
			end
		end
	end
	

endmodule
